`timescale 1ns/100ps

module eric_clapton(

    input wire [3:0] A_e, B_e, C_e,              
    input wire clk,
    input wire reset,
    output reg Yout);















endmodule
