`timescale 1ns/100ps

module mux4to1_always(f, a, sel);

	output f;
	input [3:0] a;
	input [1:0] sel;











endmodule

