`timescale 1ns/100ps

module mux2to1_primitives(f ,a, sel);

	output f;
	input [1:0] a;
	input sel;













endmodule
